`ifndef FUNCTIONS_INCLUDE_SV
    `define FUNCTIONS_INCLUDE_SV

package functions_pkg;

endpackage : functions_pkg

`endif 