// MIT License
//
// Copyright (c) 2021 Gabriele Tripi
// 
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
// -----------------------------------------------------------------------------------
// -----------------------------------------------------------------------------------
// FILE NAME : carry_lookahead_adder.sv
// DEPARTMENT : 
// AUTHOR : Gabriele Tripi
// AUTHOR'S EMAIL : tripi.gabriele2002@gmail.com
// -----------------------------------------------------------------------------------
// RELEASE HISTORY
// VERSION : 1.0 
// DATE : 28 / 10 / 2021
// DESCRIPTION : Carry Lookahead Adder, it perform binary addition in O(log(n)) time. 
//               In this file there are two modules: one for the single block and one  
//               for the entire adder (which is composed by several CLA blocks).
//               The CLA adder can take a carry as an input.
// -----------------------------------------------------------------------------------
// KEYWORDS :
// -----------------------------------------------------------------------------------
// PARAMETERS
// PARAM NAME  : RANGE   : DESCRIPTION              : DEFAULT 
// DATA_WIDTH  :    /    : I/O number of bits       : 32
// BLOCK_WIDTH :    /    : Number of bit in a block : 4
// -----------------------------------------------------------------------------------

module carry_lookahead_adder #(

  // Number of bits in a word
  parameter DATA_WIDTH = 32,

  // Number of bits computed in a CLA block
  parameter BLOCK_WIDTH = 4
) 
(
  input  logic [DATA_WIDTH - 1:0] operand_A_i,
  input  logic [DATA_WIDTH - 1:0] operand_B_i,
  input  logic                    carry_i,

  output logic [DATA_WIDTH - 1:0] result_o,
  output logic                    carry_o
);

//------------//
// PARAMETERS //
//------------//

  // Total number of CLA block 
  localparam CLA_BLOCKS = DATA_WIDTH / BLOCK_WIDTH;

//------------//
//  DATAPATH  //
//------------//

  // Carry input / output of every CLA block
  logic [CLA_BLOCKS - 1:0] cla_carry;

  genvar i;
  generate

    for (i = 0; i < CLA_BLOCKS; i++) begin 
      CLA_block N_th_CLA_block (
        .cla_operand_A_i (operand_A_i[(BLOCK_WIDTH * i) +: BLOCK_WIDTH]),
        .cla_operand_B_i (operand_B_i[(BLOCK_WIDTH * i) +: BLOCK_WIDTH]),
        .cla_carry_i     ((i == 0) ? carry_i : cla_carry[i - 1]        ),
        .cla_result_o    (result_o[(BLOCK_WIDTH * i) +: BLOCK_WIDTH]   ),
        .cla_carry_o     (cla_carry[i]                                 )
      );
    end

  endgenerate

  // Carry out is the carry generated by the last CLA block
  assign carry_o = cla_carry[CLA_BLOCKS - 1];

endmodule

module CLA_block #(

  // Number of bits computed in a CLA block
  BLOCK_WIDTH = 4
)
(
  input  logic [BLOCK_WIDTH - 1:0] cla_operand_A_i,
  input  logic [BLOCK_WIDTH - 1:0] cla_operand_B_i,
  input  logic                     cla_carry_i,

  output logic [BLOCK_WIDTH - 1:0] cla_result_o,
  output logic                     cla_carry_o
);

//------------//
// PARAMETERS //
//------------//

  // Nets inout
  localparam IN = 1;
  localparam OUT = 0;

//------------//
//  DATAPATH  //
//------------//

  // Carry bit produced by each sum bit 
  logic [IN:OUT][BLOCK_WIDTH - 1:0] carry;

  // Result of the xor between A and B
  logic [BLOCK_WIDTH - 1:0] AB_xor;

      // Ripple carry
      always_comb begin : rc_adder_logic
        for (int i = 0; i < BLOCK_WIDTH; i++) begin 
          AB_xor[i] = cla_operand_A_i[i] ^ cla_operand_B_i[i];

          // The first Full-Adder takes the external carry in
          carry[IN][i] = (i == 0) ? cla_carry_i : carry[OUT][i - 1];
          cla_result_o[i] = AB_xor[i] ^ carry[IN][i];
          carry[OUT][i] = (AB_xor[i] & carry[IN][i]) | (cla_operand_A_i[i] & cla_operand_B_i[i]);
        end
      end : rc_adder_logic

  // Generation and propagation nets
  logic [BLOCK_WIDTH - 1:0] c_generate, c_propagate;
  logic [BLOCK_WIDTH - 2:0] and_cgen, or_cgen; 

      always_comb begin : carry_logic
        for (int j = 0; j < BLOCK_WIDTH; j++) begin : generate_propagate_logic 
          c_generate[j] = cla_operand_A_i[j] & cla_operand_B_i[j]; 
          c_propagate[j] = cla_operand_A_i[j] | cla_operand_B_i[j]; 
        end : generate_propagate_logic

          // Carry generation logic
          for (int k = 0; k < BLOCK_WIDTH - 1; k++) begin : carry_gen_logic
            if (k == 0) begin 
              and_cgen[0] = c_generate[0] & c_propagate[1];
              or_cgen[0] = and_cgen[0] | c_generate[1];
            end else begin 
              and_cgen[k] = or_cgen[k - 1] & c_propagate[k + 1];
              or_cgen[k] = and_cgen[k] | c_generate[k + 1];
            end
          end : carry_gen_logic
      end : carry_logic

  assign cla_carry_o = or_cgen[BLOCK_WIDTH - 2] | (&c_propagate & cla_carry_i);

endmodule
